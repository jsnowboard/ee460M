module parkingMeterTop(CLK, UP, DWN, LEFT, RIGHT, sevenSeg);
input CLK, UP, DWN, LEFT, RIGHT;
output [3:0] sevenSeg;


endmodule
